set_property PACKAGE_PIN J15 [get_ports A]
set_property IOSTANDARD LVCMOS33 [get_ports A]
set_property PACKAGE_PIN L16 [get_ports B]
set_property IOSTANDARD LVCMOS33 [get_ports B]
set_property PACKAGE_PIN H17 [get_ports F_AND]
set_property PACKAGE_PIN K15 [get_ports F_NOT]
set_property PACKAGE_PIN J13 [get_ports F_OR]
set_property IOSTANDARD LVCMOS33 [get_ports F_AND]
set_property IOSTANDARD LVCMOS33 [get_ports F_NOT]
set_property IOSTANDARD LVCMOS33 [get_ports F_OR]
